package adder_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "item.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "sb.sv"
  `include "agent.sv"
  `include "env.sv"
  `include "sequence.sv"
  `include "test.sv"
endpackage : adder_pkg
