interface adder_if();
  logic [31:0] sum_in1;
  logic [31:0] sum_in2;
  logic [31:0] sum_out;
  logic carry_bit_out;
endinterface
